module serial()

endmodule
